// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// simmem

// This modules assumes that no capacity overflow occurs.

module simmem_delay_banks #(
  // Width of the messages, including identifier
)(

);

  // To be implemented, similarly to the delay bank

endmodule
